module video_tb ();

    // Test video playback on the main top level module



    


endmodule