// This is the controller used to initialize first load up of data into buffers before the data_FSM takes over for the rest of the operations



module startup_FSM (

);















endmodule