module vieo_playbak (

);
    // VGA controller




    // Bank counter



    // Counters

endmodule