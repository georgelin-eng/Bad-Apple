module BRAM_tb()
    

endmodule