// Testing environment so see that all the clock enable signals have the right frequency and are only high
// for a single clock cycle




