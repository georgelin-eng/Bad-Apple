///////////////////////////////////
// Buffer size: 1s audio (256kb) //
///////////////////////////////////

